module cache_sel
(
    
)